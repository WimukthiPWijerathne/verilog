module fulladder(
    inpput wire a,
    input wire b,
    input wire cin,
    output wire cout,
    output wire sum
);

    assgin {cout, sum} = a + b + cin;



    endmodule
    